module lab05part01();
endmodule
