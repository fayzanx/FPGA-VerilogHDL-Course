module lab05part02(
    output [6:0]HEX3, HEX2, HEX1, HEX0,
    input  [9:0]SW
);



endmodule
