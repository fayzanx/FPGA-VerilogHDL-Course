module main(input X,Y, output A, B);
	base_halfAdder(1'b1, 1'b1, A, B);
endmodule